module blok_ron (c,wreg,
d_bus, ax,ay,x,y, int_save, int_load);
input c,wreg, int_save, int_load ;
input [7:0] d_bus;
input [3:0] ax, ay;
output [7:0] x,y;
 reg [7:0] x,y;
reg [7:0] ron [3:0]; 
reg [7:0] prev_ron [3:0]; 
 always begin 
 x=ron[ax]; y=ron[ay]; end
 always @(posedge c) 
 begin
	if (wreg)
	begin
		ron[ax] = d_bus;
		if(int_save)
		begin
			prev_ron[0] <= ron[0];
			prev_ron[1] <= ron[1];
			prev_ron[2] <= ron[2];
			prev_ron[3] <= ron[3];
			
			
			ron[0] <= 8'b0;
			ron[1] <= 8'b0;
			ron[2] <= 8'b0;
			ron[3] <= 8'b0;
		end
		else if (int_load)
		begin
			ron[0] <= prev_ron[0];
			ron[1] <= prev_ron[1];
			ron[2] <= prev_ron[2];
			ron[3] <= prev_ron[3];
		end			
	end
end

endmodule